Begin3
Language:    SV, 850, Swedish
Title:       FED
Description: En radbrytande textredigerare med f�rgmarkering av syntax och mer �n s�
Keywords:    text, redigerare
End
